library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
entity InstrMemory is
port (address : in std_logic_vector (4 downto 0);
data : out std_logic_vector (31 downto 0));
end entity InstrMemory;

architecture beh of InstrMemory is
type mem is array (0 to 31) of std_logic_vector(31 downto 0);
constant memInstr : mem := (
"00000000011100000000100000010011",
"00001111110000010000001000010111",
"11111111110000100000001000010011",
"00001111110000010000001010010111",
"00000001000000101000001010010011",
"01000000000000000000011010110111",
"11111111111101101000011010010011",
"00000010000010000000001001100011",--
"00000000000000100010010000000011",
--"01000001111101000101010010010011",
--"00000000100101000100010100110011",
--"00000000000101001111010010010011",
--"00000000100101010000010100110011",
--abs instruction
"00000000000001000001010100010011",
"00000000010000100000001000010011",
"11111111111110000000100000010011",
"00000000110101010010010110110011",
"11111110000001011000010011100011",--
"00000000000001010000011010110011",
"11111110000111111111000011101111",--
"00000000110100101010000000100011",
"00000000000000000000000011101111",--
"00000000000000000000000000010011",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000"


);
begin
data <= memInstr(to_integer(unsigned(address)));
end architecture beh;