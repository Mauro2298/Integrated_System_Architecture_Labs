LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

USE WORK.dictionary.ALL;

ENTITY RF IS
	PORT(
		RF_IN_RS1 : IN STD_LOGIC_VECTOR(NBIT_RF_ADD-1 DOWNTO 0);
		RF_IN_RS2 : IN STD_LOGIC_VECTOR(NBIT_RF_ADD-1 DOWNTO 0);
		RF_IN_RD : IN STD_LOGIC_VECTOR(NBIT_RF_ADD-1 DOWNTO 0);
		RF_IN_WR_RD : IN STD_LOGIC;
		RF_IN_RD_DT : IN STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0);
		
		RF_IN_RST : IN STD_LOGIC;
		RF_IN_CLK : IN STD_LOGIC;
		
		RF_OUT_RS1_DT : OUT STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0);
		RF_OUT_RS2_DT : OUT STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0)
	);
END ENTITY RF;

ARCHITECTURE structural OF RF IS

	COMPONENT decoder IS
		PORT(
			DEC_IN : IN STD_LOGIC_VECTOR(NBIT_RF_ADD-1 DOWNTO 0);
			DEC_OUT : OUT STD_LOGIC_VECTOR((2**NBIT_RF_ADD)-1 DOWNTO 0)
	);
	END COMPONENT;

	COMPONENT n_bit_register IS 
		generic (n_bit: INTEGER);
		port (data_in: IN STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0);
		    CLK, reset, enable: IN std_logic;
		    data_out: OUT STD_LOGIC_VECTOR(n_bit - 1 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT mux32to1 IS
	PORT(
		MUX32_IN_DT : IN DATA_BUS_32;
		MUX32_IN_SL : IN STD_LOGIC_VECTOR (NBIT_RF_ADD-1 DOWNTO 0);
		MUX32_OUT : OUT STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0)
	);
	END COMPONENT;

SIGNAL FROM_DEC, REG_EN : STD_LOGIC_VECTOR((2**NBIT_RF_ADD)-1 DOWNTO 0);

SIGNAL REG_OUT : DATA_BUS_32;

BEGIN

	

	DEC: decoder PORT MAP(
						DEC_IN => RF_IN_RD,
						DEC_OUT => FROM_DEC
				);

	RF_REGS : FOR REG_INDEX IN 0 TO (2**NBIT_RF_ADD)-1 GENERATE
	BEGIN
	
		REG_EN(REG_INDEX) <= FROM_DEC(REG_INDEX) AND RF_IN_WR_RD;

		REG: n_bit_register GENERIC MAP (n_bit => NBIT)
							PORT MAP(
									data_in => RF_IN_RD_DT,
									CLK => RF_IN_CLK,
									reset => RF_IN_RST,
									enable => REG_EN(REG_INDEX),
									data_out => REG_OUT(REG_INDEX)
							);
	
	END GENERATE RF_REGS; 

	MUX_RS1: mux32to1 PORT MAP (
						MUX32_IN_DT => REG_OUT,
						MUX32_IN_SL => RF_IN_RS1,
						MUX32_OUT => RF_OUT_RS1_DT
					);

	MUX_RS2: mux32to1 PORT MAP (
						MUX32_IN_DT => REG_OUT,
						MUX32_IN_SL => RF_IN_RS2,
						MUX32_OUT => RF_OUT_RS2_DT
					);

END structural;