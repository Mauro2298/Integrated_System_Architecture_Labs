LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

USE WORK.dictionary.ALL;

ENTITY FW_unit IS 
	PORT(
		FW_IN_RS1_EX : IN STD_LOGIC_VECTOR (NBIT_RF_ADD-1 DOWNTO 0);
		FW_IN_RS2_EX : IN STD_LOGIC_VECTOR (NBIT_RF_ADD-1 DOWNTO 0);
		FW_IN_RD_M : IN STD_LOGIC_VECTOR (NBIT_RF_ADD-1 DOWNTO 0);
		FW_IN_RD_WB : IN STD_LOGIC_VECTOR (NBIT_RF_ADD-1 DOWNTO 0);
		
		FW_IN_WB_M : IN STD_LOGIC;
		FW_IN_WB_WB : IN STD_LOGIC;
		
		FW_OUT_FW_A_M : OUT STD_LOGIC;
		FW_OUT_FW_A_WB : OUT STD_LOGIC;
		FW_OUT_FW_B_M : OUT STD_LOGIC;
		FW_OUT_FW_B_WB : OUT STD_LOGIC
	);
END ENTITY;

ARCHITECTURE behavioral OF FW_unit IS
	
BEGIN

	FW_OUT_FW_A_M <= '1' WHEN ((FW_IN_RS1_EX = FW_IN_RD_M) AND FW_IN_WB_M = '1') ELSE '0';
	
	FW_OUT_FW_A_WB <= '1' WHEN ((FW_IN_RS1_EX = FW_IN_RD_WB) AND FW_IN_WB_WB ='1') ELSE '0';

	FW_OUT_FW_B_M <= '1' WHEN ((FW_IN_RS2_EX = FW_IN_RD_M) AND FW_IN_WB_M = '1') ELSE '0';
	
	FW_OUT_FW_B_WB <= '1' WHEN ((FW_IN_RS2_EX = FW_IN_RD_WB) AND FW_IN_WB_WB = '1') ELSE '0';
		
END ARCHITECTURE behavioral;