LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY int_comparator IS
        GENERIC (N : INTEGER);
        PORT (
            INT_CMP_IN_A : IN STD_LOGIC_VECTOR (N-1 DOWNTO 0);
            INT_CMP_IN_B : IN STD_LOGIC_VECTOR (N-1 DOWNTO 0);
            INT_CMP_OUT : OUT STD_LOGIC_VECTOR (N-1 DOWNTO 0)
        );
END ENTITY;

ARCHITECTURE behavioral OF int_comparator IS

    SIGNAL RESULT : STD_LOGIC_VECTOR (N-1 DOWNTO 0);

BEGIN

    --THE COMPARE OPERATION EXPLOITS A SUBTRACTOR
    RESULT <= STD_LOGIC_VECTOR( SIGNED(INT_CMP_IN_A) - SIGNED(INT_CMP_IN_B) );

    --THE OUTPUT VALUE IS DERIVED BY THE SIGN OF THE RESULT
    INT_CMP_OUT <= STD_LOGIC_VECTOR(TO_UNSIGNED(0,N-1)) & RESULT(N-1);

END behavioral;
