LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

USE WORK.BF.ALL;

ENTITY MBE IS 
    --GENERIC (NBIT : INTEGER := 33);
    PORT(
        MBE_IN_MULTIPLICAND : IN STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0);
        MBE_IN_MULTIPLIER : IN STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0);
        MBE_OUT_RESULT : OUT STD_LOGIC_VECTOR(COLUMN_NUMBER -1 DOWNTO 0)
    );
END MBE;

ARCHITECTURE BEH OF MBE IS

	COMPONENT MBE_Multiplier IS 
		--GENERIC (NBIT : INTEGER := 33);
		PORT(
		    MBE_IN_MULTIPLICAND : IN STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0);
		    MBE_IN_MULTIPLIER : IN STD_LOGIC_VECTOR(NBIT-1 DOWNTO 0);
		    MBE_OUT_RESULT : OUT STD_LOGIC_VECTOR(COLUMN_NUMBER DOWNTO 0)
		);
	END COMPONENT;

	SIGNAL OUT_RES : STD_LOGIC_VECTOR(COLUMN_NUMBER DOWNTO 0);
BEGIN

	MBE_COMP: MBE_Multiplier PORT MAP(
        MBE_IN_MULTIPLICAND => MBE_IN_MULTIPLICAND,
        MBE_IN_MULTIPLIER => MBE_IN_MULTIPLIER,
        MBE_OUT_RESULT => OUT_RES
    );

	MBE_OUT_RESULT <= OUT_RES(COLUMN_NUMBER - 1 DOWNTO 0);
END BEH;
