library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package packa is
type stage is array (0 to 10) of std_logic_vector(12 downto 0);
end package;
