PACKAGE constants IS
	constant N : natural := 4;
END constants;
