LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.dictionary.ALL;

ENTITY immediate_gen IS
	
	PORT(
		IMM_GEN_IN_INST : IN STD_LOGIC_VECTOR (NBIT_INST-1 DOWNTO 0);
		IMM_GEN_OUT_IMM : OUT STD_LOGIC_VECTOR (NBIT_INST-1 DOWNTO 0)
	);

END ENTITY immediate_gen;

ARCHITECTURE behavioral OF immediate_gen IS

SIGNAL SIGN_EXT : STD_LOGIC_VECTOR(26 DOWNTO 0);

BEGIN

SIGN_EXT <= (OTHERS=>IMM_GEN_IN_INST(31));

	IMM_GEN_OUT_IMM <= 
						IMM_GEN_IN_INST(31 DOWNTO 12) & STD_LOGIC_VECTOR(TO_UNSIGNED(0,12))
						WHEN ( IMM_GEN_IN_INST(NBIT_OPCODE-1 DOWNTO 0) = LUI ) OR ( IMM_GEN_IN_INST(NBIT_OPCODE-1 DOWNTO 0) = AUIPC ) ELSE
						
						SIGN_EXT(19 DOWNTO 0) & IMM_GEN_IN_INST(31 DOWNTO 20) 
						WHEN ( IMM_GEN_IN_INST(NBIT_OPCODE-1 DOWNTO 0) = IMMA ) OR ( IMM_GEN_IN_INST(NBIT_OPCODE-1 DOWNTO 0) = IMML ) ELSE
						
						SIGN_EXT(19 DOWNTO 0) & IMM_GEN_IN_INST(31 DOWNTO 25) & IMM_GEN_IN_INST(11 DOWNTO 7) 
						WHEN ( IMM_GEN_IN_INST(NBIT_OPCODE-1 DOWNTO 0) = S ) ELSE
						
						SIGN_EXT(10 DOWNTO 0) & IMM_GEN_IN_INST(31) & IMM_GEN_IN_INST(19 DOWNTO 12) & IMM_GEN_IN_INST(20) & IMM_GEN_IN_INST(30 DOWNTO 21) & '0'
						WHEN ( IMM_GEN_IN_INST(NBIT_OPCODE-1 DOWNTO 0) = J ) ELSE
						
						SIGN_EXT(18 DOWNTO 0) & IMM_GEN_IN_INST(31) & IMM_GEN_IN_INST(7) & IMM_GEN_IN_INST(30 DOWNTO 25) & IMM_GEN_IN_INST(11 DOWNTO 8) & '0'
						WHEN ( IMM_GEN_IN_INST(NBIT_OPCODE-1 DOWNTO 0) = B ) ELSE
						
						STD_LOGIC_VECTOR(TO_UNSIGNED(0,27)) & IMM_GEN_IN_INST(24 DOWNTO 20) 
						WHEN ( IMM_GEN_IN_INST(NBIT_OPCODE-1 DOWNTO 0) = IMMS ) ELSE 
						
						(OTHERS=>'0');

END ARCHITECTURE behavioral;