library verilog;
use verilog.vl_types.all;
entity tb_RISCV is
end tb_RISCV;
