LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

USE WORK.dictionary.ALL;

ENTITY CTRL_unit IS
	PORT(
		CTRL_IN_OPCODE : IN STD_LOGIC_VECTOR(NBIT_OPCODE-1 DOWNTO 0);
		
		CTRL_OUT_IMML : OUT STD_LOGIC;
		CTRL_OUT_IMMA : OUT STD_LOGIC;
		CTRL_OUT_IMMS : OUT STD_LOGIC;
		CTRL_OUT_B : OUT STD_LOGIC;
		CTRL_OUT_J : OUT STD_LOGIC;
		CTRL_OUT_LUI : OUT STD_LOGIC;
		CTRL_OUT_AUIPC : OUT STD_LOGIC;
		CTRL_OUT_S : OUT STD_LOGIC;
		CTRL_OUT_RA : OUT STD_LOGIC;
		
		CTRL_OUT_EX : OUT STD_LOGIC;
		CTRL_OUT_WB : OUT STD_LOGIC
	);
END ENTITY;

ARCHITECTURE behavioral OF CTRL_unit IS

BEGIN

	CTRL_OUT_IMML <= '1' WHEN CTRL_IN_OPCODE = IMML ELSE '0';
	CTRL_OUT_IMMA <= '1' WHEN CTRL_IN_OPCODE = IMMA ELSE '0';
	CTRL_OUT_IMMS <= '1' WHEN CTRL_IN_OPCODE = IMMS ELSE '0';
	CTRL_OUT_B <= '1' WHEN CTRL_IN_OPCODE = B ELSE '0';
	CTRL_OUT_J <= '1' WHEN CTRL_IN_OPCODE = J ELSE '0';
	CTRL_OUT_LUI <= '1' WHEN CTRL_IN_OPCODE = LUI ELSE '0';
	CTRL_OUT_AUIPC <= '1' WHEN CTRL_IN_OPCODE = AUIPC ELSE '0';
	CTRL_OUT_S <= '1' WHEN CTRL_IN_OPCODE = S ELSE '0';
	CTRL_OUT_RA <= '1' WHEN CTRL_IN_OPCODE = RA ELSE '0';

	CTRL_OUT_EX <= '1' WHEN ( (CTRL_IN_OPCODE = IMML) OR (CTRL_IN_OPCODE = IMMA) OR (CTRL_IN_OPCODE = IMMS) OR (CTRL_IN_OPCODE = RA) OR (CTRL_IN_OPCODE = S) OR (CTRL_IN_OPCODE = AUIPC) OR (CTRL_IN_OPCODE = B) ) ELSE '0';
	
	CTRL_OUT_WB <= '1' WHEN ( (CTRL_IN_OPCODE = IMML) OR (CTRL_IN_OPCODE = IMMA) OR (CTRL_IN_OPCODE = IMMS) OR (CTRL_IN_OPCODE = RA) OR (CTRL_IN_OPCODE = AUIPC) OR (CTRL_IN_OPCODE = LUI) OR (CTRL_IN_OPCODE = J) ) ELSE '0';

END ARCHITECTURE behavioral;